Output Before Switching
V1 1 0 dc 1V
R1 X 1 1
C1 X 0 1u ic=0
R2 X 3 2
V2 3 0 dc 2V
.tran 10p 10u uic

.control
run
set gnuplot_terminal=png/quit
gnuplot ../figs/2_7 v(X)
.endc

.end
