Output After Switching
R1 X 0 1
C1 X 0 1u ic=1.33
R2 X 3 2
V2 3 0 dc 2V
.tran 10p 10u uic

.control
run
set gnuplot_terminal=png/quit
gnuplot ../figs/3_5 v(X) 
.endc

.end
